
//--xuezhen--

`include "defines.v"

module SimTop(
    input         clock,
    input         reset,

    input  [63:0] io_logCtrl_log_begin,
    input  [63:0] io_logCtrl_log_end,
    input  [63:0] io_logCtrl_log_level,
    input         io_perfInfo_clean,
    input         io_perfInfo_dump,

    output        io_uart_out_valid,
    output [7:0]  io_uart_out_ch,
    output        io_uart_in_valid,
    input  [7:0]  io_uart_in_ch
);

// if_stage
wire [63 : 0] pc;
wire [31 : 0] inst;
wire inst_ena;

// id_stage
// id_stage -> regfile
wire rs1_r_ena;
wire [4 : 0]rs1_r_addr;
wire rs2_r_ena;
wire [4 : 0]rs2_r_addr;
wire rd_w_ena;
wire [4 : 0]rd_w_addr;
// id_stage -> exe_stage
wire [4 : 0]inst_type;
wire [7 : 0]inst_opcode;
wire [`REG_BUS]op1;
wire [`REG_BUS]op2;
wire [2:0] alumem_reg;

// id_stage -> if_stage
wire [1  : 0]mpc;
wire [63 : 0]imm;
wire [2  : 0]jump;

//id_stage -> mem_stage
wire wen;
wire[63 : 0] wdata;
wire[63 : 0] wmask;
// regfile -> id_stage
wire [`REG_BUS] r_data1;
wire [`REG_BUS] r_data2;
// regfile -> difftest
wire [`REG_BUS] regs[0 : 31];

// exe_stage
// exe_stage -> other stage
wire [4 : 0]inst_type_o;
wire [`REG_BUS]memr_data;
wire [`REG_BUS]exe_data;
wire zero;
// exe_stage -> regfile
wire [`REG_BUS]rd_data;


// Access memory
reg [63:0] rdata;
reg [63:0] rdata2;
RAMHelper RAMHelper(
  .clk              (clock),
  .en               (1),
  .rIdx             ((pc - `PC_START) >> 3),
  .rdata            (rdata),
  .wIdx             ((exe_data - `PC_START) >> 3),
  .wdata            (wdata),
  .wmask            (wmask),
  .wen              (wen)
);
assign inst = pc[2] ? rdata[63 : 32] : rdata[31 : 0];


RAMHelper RAMHelperdata(
  .clk              (clock),
  .en               (1),
  .rIdx             ((exe_data - `PC_START) >> 3),
  .rdata            (rdata2),
  .wIdx             (0),
  .wdata            (0),
  .wmask            (0),
  .wen              (0)
);
assign memr_data = rdata2;
//exe_data[2] ? rdata2[63 : 32] : rdata2[31 : 0];

if_stage If_stage(
  .clk(clock),
  .rst(reset),
 // .mpc(mpc),
  .imm(imm),
  .jump(jump),
  .pc_o(pc),
  .zero(zero),
  .r_data1         (r_data1)
);

id_stage Id_stage(
  .rst              (reset),
  .inst             (inst),
  .rs1_data         (r_data1),
  .rs2_data         (r_data2),
  .inst_addr        (pc),
  .exe_data(exe_data),
  
  .rs1_r_ena        (rs1_r_ena),
  .rs1_r_addr       (rs1_r_addr),
  .rs2_r_ena        (rs2_r_ena),
  .rs2_r_addr       (rs2_r_addr),
  .rd_w_ena         (rd_w_ena),
  .rd_w_addr        (rd_w_addr),
  .inst_type        (inst_type),
  .inst_opcode      (inst_opcode),
  .op1              (op1),
  .op2              (op2),
  .mpc              (mpc),
  .imm              (imm),
  .jump_o           (jump),
  .alumem_reg(alumem_reg),
  
  .mem_wen(wen),       // Mem write
  .mem_wdata(wdata),
  .wmask            (wmask)
);

exe_stage Exe_stage(
  .rst              (reset),
  .inst_type_i      (inst_type),
  .inst_opcode      (inst_opcode),
  .op1              (op1),
  .op2              (op2),
  .inst             (inst),
  .alumem_reg(alumem_reg),
  .memr_data(memr_data),
  .exe_data(exe_data),
  .inst_type_o      (inst_type_o),
  .rd_data          (rd_data),
  .zero(zero)
);

regfile Regfile(
  .clk              (clock),
  .rst              (reset),
  .w_addr           (rd_w_addr),
  .w_data           (rd_data),
  .w_ena            (rd_w_ena),
  
  .r_addr1          (rs1_r_addr),
  .r_data1          (r_data1),
  .r_ena1           (rs1_r_ena),
  .r_addr2          (rs2_r_addr),
  .r_data2          (r_data2),
  .r_ena2           (rs2_r_ena),

  .regs_o           (regs)
);


// Difftest
reg cmt_wen;
reg [7:0]cmt_wdest;
reg [`REG_BUS] cmt_wdata;
reg [`REG_BUS] cmt_pc;
reg [31:0]cmt_inst;
reg vaild;
reg skip;
reg [63:0] cycleCnt;
reg [63:0] instrCnt;

always @(posedge clock) begin
  if (reset) begin
    {cmt_wen, cmt_wdest, cmt_wdata, cmt_pc, cmt_inst, vaild, cycleCnt, instrCnt} = 0;
  end
  else begin
    cmt_wen = rd_w_ena;
    cmt_wdest = {3'd0, rd_w_addr};
    cmt_wdata = rd_data;
    cmt_pc = pc;
    cmt_inst = inst;
    vaild = 1'd1;

    // Skip comparison of the first instruction
    // Because the result required to commit cannot be calculated in time before first InstrCommit during verilator simulation
    // Maybe you can avoid it in pipeline
    skip = pc == `PC_START;
    
    cycleCnt += 1;
    instrCnt += 1;
  end
end

DifftestInstrCommit DifftestInstrCommit(
  .clock              (clock),
  .coreid             (0),
  .index              (0),
  .valid              (vaild),
  .pc                 (cmt_pc),
  .instr              (cmt_inst),
  .skip               (skip),
  .isRVC              (0),
  .scFailed           (0),
  .wen                (cmt_wen),
  .wdest              (cmt_wdest),
  .wdata              (cmt_wdata)
);

DifftestArchIntRegState DifftestArchIntRegState (
  .clock              (clock),
  .coreid             (0),
  .gpr_0              (regs[0]),
  .gpr_1              (regs[1]),
  .gpr_2              (regs[2]),
  .gpr_3              (regs[3]),
  .gpr_4              (regs[4]),
  .gpr_5              (regs[5]),
  .gpr_6              (regs[6]),
  .gpr_7              (regs[7]),
  .gpr_8              (regs[8]),
  .gpr_9              (regs[9]),
  .gpr_10             (regs[10]),
  .gpr_11             (regs[11]),
  .gpr_12             (regs[12]),
  .gpr_13             (regs[13]),
  .gpr_14             (regs[14]),
  .gpr_15             (regs[15]),
  .gpr_16             (regs[16]),
  .gpr_17             (regs[17]),
  .gpr_18             (regs[18]),
  .gpr_19             (regs[19]),
  .gpr_20             (regs[20]),
  .gpr_21             (regs[21]),
  .gpr_22             (regs[22]),
  .gpr_23             (regs[23]),
  .gpr_24             (regs[24]),
  .gpr_25             (regs[25]),
  .gpr_26             (regs[26]),
  .gpr_27             (regs[27]),
  .gpr_28             (regs[28]),
  .gpr_29             (regs[29]),
  .gpr_30             (regs[30]),
  .gpr_31             (regs[31])
);

DifftestTrapEvent DifftestTrapEvent(
  .clock              (clock),
  .coreid             (0),
  .valid              (inst[6:0] == 7'h6b),
  .code               (regs[10][7:0]),
  .pc                 (cmt_pc),
  .cycleCnt           (cycleCnt),
  .instrCnt           (instrCnt)
);

DifftestCSRState DifftestCSRState(
  .clock              (clock),
  .coreid             (0),
  .priviledgeMode     (0),
  .mstatus            (0),
  .sstatus            (0),
  .mepc               (0),
  .sepc               (0),
  .mtval              (0),
  .stval              (0),
  .mtvec              (0),
  .stvec              (0),
  .mcause             (0),
  .scause             (0),
  .satp               (0),
  .mip                (0),
  .mie                (0),
  .mscratch           (0),
  .sscratch           (0),
  .mideleg            (0),
  .medeleg            (0)
);

DifftestArchFpRegState DifftestArchFpRegState(
  .clock              (clock),
  .coreid             (0),
  .fpr_0              (0),
  .fpr_1              (0),
  .fpr_2              (0),
  .fpr_3              (0),
  .fpr_4              (0),
  .fpr_5              (0),
  .fpr_6              (0),
  .fpr_7              (0),
  .fpr_8              (0),
  .fpr_9              (0),
  .fpr_10             (0),
  .fpr_11             (0),
  .fpr_12             (0),
  .fpr_13             (0),
  .fpr_14             (0),
  .fpr_15             (0),
  .fpr_16             (0),
  .fpr_17             (0),
  .fpr_18             (0),
  .fpr_19             (0),
  .fpr_20             (0),
  .fpr_21             (0),
  .fpr_22             (0),
  .fpr_23             (0),
  .fpr_24             (0),
  .fpr_25             (0),
  .fpr_26             (0),
  .fpr_27             (0),
  .fpr_28             (0),
  .fpr_29             (0),
  .fpr_30             (0),
  .fpr_31             (0)
);

endmodule
